//Convert signal from TIA to VGA buffer

//Notes: Image is scanlines 40-231, Pixels 68-227

module VGA(input  logic [8:0]  ScanLine,
			  input  logic [7:0]  xPos);
			  input logic [6:0]  CurColor

endmodule

//Top-level module for 2600

module a2600();
endmodule
